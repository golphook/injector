module main

//const target_name = "dummy_prog.exe"
const target_name = "csgo.exe"
const to_clear = [".rsrc", ".reloc", ".00cfg"]
//const dll_ressource = 'ressources/cool_dll.dll'
const dll_ressource = "ressources/golphook.dll"
