module main

const target_name = "csgo.exe"
