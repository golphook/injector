module main

const target_name = "csgo.exe"
const to_clear = [".rsrc", ".reloc", ".00cfg"]
