module main

const target_name = "csgo.exe"
const to_clear = [".rsrc", ".reloc", ".00cfg"]

const latest_version = "to_rep_ci"
